`timescale 1ns / 1ps

module eth_crc32(
	input clk,
	input en,
	input rst,
	input [7:0]dat,
	output [31:0]crc
	);

reg [31:0]c = 32'hFFFFFFFF;
reg [31:0]nxt;

wire [7:0]d = { dat[0],dat[1],dat[2],dat[3],dat[4],dat[5],dat[6],dat[7] };

assign crc = {
	c[0],c[1],c[2],c[3],c[4],c[5],c[6],c[7],
	c[8],c[9],c[10],c[11],c[12],c[13],c[14],c[15],
	c[16],c[17],c[18],c[19],c[20],c[21],c[22],c[23],
	c[24],c[25],c[26],c[27],c[28],c[29],c[30],c[31]
	};

always_comb begin 
	nxt[0] = c[24]^c[30]^d[0]^d[6];
	nxt[1] = c[24]^c[25]^c[30]^c[31]^d[0]^d[1]^d[6]^d[7];
	nxt[2] = c[24]^c[25]^c[26]^c[30]^c[31]^d[0]^d[1]^d[2]^d[6]^d[7];
	nxt[3] = c[25]^c[26]^c[27]^c[31]^d[1]^d[2]^d[3]^d[7];
	nxt[4] = c[24]^c[26]^c[27]^c[28]^c[30]^d[0]^d[2]^d[3]^d[4]^d[6];
	nxt[5] = c[24]^c[25]^c[27]^c[28]^c[29]^c[30]^c[31]^d[0]^d[1]^d[3]^d[4]^d[5]^d[6]^d[7];
	nxt[6] = c[25]^c[26]^c[28]^c[29]^c[30]^c[31]^d[1]^d[2]^d[4]^d[5]^d[6]^d[7];
	nxt[7] = c[24]^c[26]^c[27]^c[29]^c[31]^d[0]^d[2]^d[3]^d[5]^d[7];
	nxt[8] = c[0]^c[24]^c[25]^c[27]^c[28]^d[0]^d[1]^d[3]^d[4];
	nxt[9] = c[1]^c[25]^c[26]^c[28]^c[29]^d[1]^d[2]^d[4]^d[5];
	nxt[10] = c[2]^c[24]^c[26]^c[27]^c[29]^d[0]^d[2]^d[3]^d[5];
	nxt[11] = c[3]^c[24]^c[25]^c[27]^c[28]^d[0]^d[1]^d[3]^d[4];
	nxt[12] = c[4]^c[24]^c[25]^c[26]^c[28]^c[29]^c[30]^d[0]^d[1]^d[2]^d[4]^d[5]^d[6];
	nxt[13] = c[5]^c[25]^c[26]^c[27]^c[29]^c[30]^c[31]^d[1]^d[2]^d[3]^d[5]^d[6]^d[7];
	nxt[14] = c[6]^c[26]^c[27]^c[28]^c[30]^c[31]^d[2]^d[3]^d[4]^d[6]^d[7];
	nxt[15] = c[7]^c[27]^c[28]^c[29]^c[31]^d[3]^d[4]^d[5]^d[7];
	nxt[16] = c[8]^c[24]^c[28]^c[29]^d[0]^d[4]^d[5];
	nxt[17] = c[9]^c[25]^c[29]^c[30]^d[1]^d[5]^d[6];
	nxt[18] = c[10]^c[26]^c[30]^c[31]^d[2]^d[6]^d[7];
	nxt[19] = c[11]^c[27]^c[31]^d[3]^d[7];
	nxt[20] = c[12]^c[28]^d[4];
	nxt[21] = c[13]^c[29]^d[5];
	nxt[22] = c[14]^c[24]^d[0];
	nxt[23] = c[15]^c[24]^c[25]^c[30]^d[0]^d[1]^d[6];
	nxt[24] = c[16]^c[25]^c[26]^c[31]^d[1]^d[2]^d[7];
	nxt[25] = c[17]^c[26]^c[27]^d[2]^d[3];
	nxt[26] = c[18]^c[24]^c[27]^c[28]^c[30]^d[0]^d[3]^d[4]^d[6];
	nxt[27] = c[19]^c[25]^c[28]^c[29]^c[31]^d[1]^d[4]^d[5]^d[7];
	nxt[28] = c[20]^c[26]^c[29]^c[30]^d[2]^d[5]^d[6];
	nxt[29] = c[21]^c[27]^c[30]^c[31]^d[3]^d[6]^d[7];
	nxt[30] = c[22]^c[28]^c[31]^d[4]^d[7];
	nxt[31] = c[23]^c[29]^d[5];
end

always @(posedge clk) begin
	if (rst) begin
		c <= 32'hFFFFFFFF;
	end else if (en) begin
		c <= nxt;
	end
end

endmodule
