
`timescale 1ns/1ps

module axi4_sram_ip #(
	parameter integer C_S00_AXI_ID_WIDTH	= 1,
	parameter integer C_S00_AXI_DATA_WIDTH	= 32,
	parameter integer C_S00_AXI_ADDR_WIDTH	= 32
	) (
	input wire  s00_axi_aclk,
	input wire  s00_axi_aresetn,
	input wire [C_S00_AXI_ID_WIDTH-1 : 0] s00_axi_awid,
	input wire [C_S00_AXI_ADDR_WIDTH-1 : 0] s00_axi_awaddr,
	input wire [7 : 0] s00_axi_awlen,
	input wire [2 : 0] s00_axi_awsize,
	input wire [1 : 0] s00_axi_awburst,
	input wire  s00_axi_awlock,
	input wire [3 : 0] s00_axi_awcache,
	input wire [2 : 0] s00_axi_awprot,
	input wire [3 : 0] s00_axi_awqos,
	input wire [3 : 0] s00_axi_awregion,
	input wire  s00_axi_awvalid,
	output wire  s00_axi_awready,
	input wire [C_S00_AXI_DATA_WIDTH-1 : 0] s00_axi_wdata,
	input wire [(C_S00_AXI_DATA_WIDTH/8)-1 : 0] s00_axi_wstrb,
	input wire  s00_axi_wlast,
	input wire  s00_axi_wvalid,
	output wire  s00_axi_wready,
	output wire [C_S00_AXI_ID_WIDTH-1 : 0] s00_axi_bid,
	output wire [1 : 0] s00_axi_bresp,
	output wire  s00_axi_bvalid,
	input wire  s00_axi_bready,
	input wire [C_S00_AXI_ID_WIDTH-1 : 0] s00_axi_arid,
	input wire [C_S00_AXI_ADDR_WIDTH-1 : 0] s00_axi_araddr,
	input wire [7 : 0] s00_axi_arlen,
	input wire [2 : 0] s00_axi_arsize,
	input wire [1 : 0] s00_axi_arburst,
	input wire  s00_axi_arlock,
	input wire [3 : 0] s00_axi_arcache,
	input wire [2 : 0] s00_axi_arprot,
	input wire [3 : 0] s00_axi_arqos,
	input wire [3 : 0] s00_axi_arregion,
	input wire  s00_axi_arvalid,
	output wire  s00_axi_arready,
	output wire [C_S00_AXI_ID_WIDTH-1 : 0] s00_axi_rid,
	output wire [C_S00_AXI_DATA_WIDTH-1 : 0] s00_axi_rdata,
	output wire [1 : 0] s00_axi_rresp,
	output wire  s00_axi_rlast,
	output wire  s00_axi_rvalid,
	input wire  s00_axi_rready
	);

axi4_sram_impl #(
	.AWIDTH(C_S00_AXI_ADDR_WIDTH),
	.DWIDTH(C_S00_AXI_DATA_WIDTH),
	.IWIDTH(C_S00_AXI_ID_WIDTH)
	) impl (
        .s00_axi_aclk(s00_axi_aclk),
        .s00_axi_aresetn(s00_axi_aresetn),
        .s00_axi_awid(s00_axi_awid),
        .s00_axi_awaddr(s00_axi_awaddr),
        .s00_axi_awlen(s00_axi_awlen),
        .s00_axi_awsize(s00_axi_awsize),
        .s00_axi_awburst(s00_axi_awburst),
        .s00_axi_awlock(s00_axi_awlock),
        .s00_axi_awcache(s00_axi_awcache),
        .s00_axi_awprot(s00_axi_awprot),
        .s00_axi_awqos(s00_axi_awqos),
        .s00_axi_awregion(s00_axi_awregion),
        .s00_axi_awvalid(s00_axi_awvalid),
        .s00_axi_awready(s00_axi_awready),
        .s00_axi_wdata(s00_axi_wdata),
        .s00_axi_wstrb(s00_axi_wstrb),
        .s00_axi_wlast(s00_axi_wlast),
        .s00_axi_wvalid(s00_axi_wvalid),
        .s00_axi_wready(s00_axi_wready),
        .s00_axi_bid(s00_axi_bid),
        .s00_axi_bresp(s00_axi_bresp),
        .s00_axi_bvalid(s00_axi_bvalid),
        .s00_axi_bready(s00_axi_bready),
        .s00_axi_arid(s00_axi_arid),
        .s00_axi_araddr(s00_axi_araddr),
        .s00_axi_arlen(s00_axi_arlen),
        .s00_axi_arsize(s00_axi_arsize),
        .s00_axi_arburst(s00_axi_arburst),
        .s00_axi_arlock(s00_axi_arlock),
        .s00_axi_arcache(s00_axi_arcache),
        .s00_axi_arprot(s00_axi_arprot),
        .s00_axi_arqos(s00_axi_arqos),
        .s00_axi_arregion(s00_axi_arregion),
        .s00_axi_arvalid(s00_axi_arvalid),
        .s00_axi_arready(s00_axi_arready),
        .s00_axi_rid(s00_axi_rid),
        .s00_axi_rdata(s00_axi_rdata),
        .s00_axi_rresp(s00_axi_rresp),
        .s00_axi_rlast(s00_axi_rlast),
        .s00_axi_rvalid(s00_axi_rvalid),
        .s00_axi_rready(s00_axi_rready)
	);

endmodule
